library verilog;
use verilog.vl_types.all;
entity lc3Pkg is
end lc3Pkg;
