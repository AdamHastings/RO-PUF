library verilog;
use verilog.vl_types.all;
entity lc3_control_sv_unit is
end lc3_control_sv_unit;
