library verilog;
use verilog.vl_types.all;
entity TransactionPkg is
end TransactionPkg;
