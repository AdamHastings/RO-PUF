library verilog;
use verilog.vl_types.all;
entity lc3_testbench is
end lc3_testbench;
