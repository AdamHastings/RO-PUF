library verilog;
use verilog.vl_types.all;
entity tb_pkg is
end tb_pkg;
