library verilog;
use verilog.vl_types.all;
entity Alu_RISC_v_unit is
end Alu_RISC_v_unit;
