package TbEnvPkg;
`include "opcodes_include.v"
parameter HALT=4'b1111;   
`include "Generator.sv"
`include "Agent.sv"
`include "ScoreBoard.sv"
`include "Driver.sv"   
`include "Environment.sv"

endpackage // TbEnvPkg
   


   