library verilog;
use verilog.vl_types.all;
entity test is
    generic(
        ADDRESS_WIDTH   : integer := 8
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of ADDRESS_WIDTH : constant is 1;
end test;
