library verilog;
use verilog.vl_types.all;
entity mem_if is
    port(
        clk             : in     vl_logic
    );
end mem_if;
