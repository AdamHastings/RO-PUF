library verilog;
use verilog.vl_types.all;
entity TbEnvPkg is
end TbEnvPkg;
