library verilog;
use verilog.vl_types.all;
entity tb_pkg_sv_unit is
end tb_pkg_sv_unit;
