library verilog;
use verilog.vl_types.all;
entity arb_if is
end arb_if;
