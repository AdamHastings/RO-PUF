package tb_pkg;
   
class Transaction;
   rand bit req;
   rand bit en;

   /*constraint creq_dist {
      req dist { 0 :/ 30, 1 :/ 70};
   }
   
   constraint cen_dist { 
      en dist { 0 :/ 5, 1 :/95 };
   }*/
   
endclass // Transaction
   
endpackage