library verilog;
use verilog.vl_types.all;
entity sram_if is
end sram_if;
