library verilog;
use verilog.vl_types.all;
entity SPM_IF is
    port(
        clk             : in     vl_logic
    );
end SPM_IF;
